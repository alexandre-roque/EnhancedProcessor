library verilog;
use verilog.vl_types.all;
entity simula is
end simula;
